package Counter24;

interface 

endpackage
package Counter;

interface 

endpackage